
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package utility is
type speed_t is (quarter, half, normal, doble);
type nbits_t is (fivebits,sixbits,sevenbits,eightbits);
end package;
 
package body utility is

end package body utility;
